/* trial module */
/* 1 inputs NOT */

module TRIAL_NOT1(
  input  IN  ,  //  input
  output O      //  output
);

//-----
// NOT 
//-----
  
  assign O = ~IN;
  
endmodule
